CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 10
2 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
170 176 283 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 148 211 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89884e-315 0
0
7 Pulser~
4 112 337 0 10 12
0 18 19 15 20 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
391 0 0
2
5.89884e-315 5.39824e-315
0
2 +V
167 171 147 0 1 3
0 17
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89884e-315 5.39306e-315
0
6 74LS48
188 888 257 0 14 29
0 9 10 11 12 21 22 2 3 4
5 6 7 8 23
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3421 0 0
2
5.89884e-315 5.38788e-315
0
6 74112~
219 329 253 0 7 32
0 17 16 15 16 17 24 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
8157 0 0
2
5.89884e-315 5.37752e-315
0
6 74112~
219 435 253 0 7 32
0 17 12 15 12 17 25 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
5572 0 0
2
5.89884e-315 5.36716e-315
0
6 74112~
219 548 252 0 7 32
0 17 14 15 14 17 26 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
5.89884e-315 5.3568e-315
0
6 74112~
219 721 246 0 7 32
0 17 13 15 13 17 27 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7361 0 0
2
5.89884e-315 5.34643e-315
0
9 2-In AND~
219 430 74 0 3 22
0 12 11 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
5.89884e-315 5.32571e-315
0
9 2-In AND~
219 586 82 0 3 22
0 14 10 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
5.89884e-315 5.30499e-315
0
9 CC 7-Seg~
183 1162 191 0 18 19
10 8 7 6 5 4 3 2 28 29
1 1 1 0 0 1 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
5.89884e-315 5.26354e-315
0
37
0 7 0 0 0 0 0 0 5 25 0 2
367 217
353 217
7 7 2 0 0 12416 0 4 11 0 0 5
920 221
1013 221
1013 294
1177 294
1177 227
8 6 3 0 0 12416 0 4 11 0 0 5
920 230
1018 230
1018 289
1171 289
1171 227
9 5 4 0 0 12416 0 4 11 0 0 5
920 239
1023 239
1023 284
1165 284
1165 227
10 4 5 0 0 12416 0 4 11 0 0 5
920 248
1028 248
1028 279
1159 279
1159 227
11 3 6 0 0 12416 0 4 11 0 0 5
920 257
1033 257
1033 269
1153 269
1153 227
12 2 7 0 0 4224 0 4 11 0 0 3
920 266
1147 266
1147 227
13 1 8 0 0 4224 0 4 11 0 0 3
920 275
1141 275
1141 227
7 1 9 0 0 4224 0 8 4 0 0 4
745 210
843 210
843 221
856 221
0 2 10 0 0 12416 0 0 4 14 0 6
579 206
600 206
600 269
838 269
838 230
856 230
0 3 11 0 0 4224 0 0 4 18 0 4
473 265
843 265
843 239
856 239
0 4 13 0 0 4096 0 0 8 13 0 3
606 117
606 228
697 228
3 2 13 0 0 8320 0 10 8 0 0 4
607 82
606 82
606 210
697 210
2 7 10 0 0 0 0 10 7 0 0 6
562 91
552 91
552 181
579 181
579 216
572 216
0 4 14 0 0 4224 0 0 7 17 0 3
469 74
469 234
524 234
0 1 14 0 0 0 0 0 10 17 0 3
505 74
505 73
562 73
3 2 14 0 0 0 0 9 7 0 0 4
451 74
506 74
506 216
524 216
2 7 11 0 0 0 0 9 6 0 0 6
406 83
396 83
396 270
473 270
473 217
459 217
1 0 12 0 0 0 0 9 0 0 25 3
406 65
375 65
375 217
3 0 15 0 0 8192 0 8 0 0 23 3
691 219
610 219
610 371
3 0 15 0 0 0 0 7 0 0 23 3
518 225
510 225
510 371
3 0 15 0 0 0 0 6 0 0 23 3
405 226
401 226
401 371
0 0 15 0 0 8336 0 0 0 26 0 3
291 326
291 371
730 371
0 4 12 0 0 0 0 0 6 25 0 3
383 217
383 235
411 235
4 2 12 0 0 0 0 4 6 0 0 6
856 248
848 248
848 177
367 177
367 217
411 217
3 3 15 0 0 0 0 2 5 0 0 4
136 328
291 328
291 226
299 226
0 4 16 0 0 8192 0 0 5 28 0 3
184 217
184 235
305 235
1 2 16 0 0 8320 0 1 5 0 0 3
160 211
160 217
305 217
5 0 17 0 0 4096 0 5 0 0 37 2
329 265
329 296
5 0 17 0 0 8192 0 8 0 0 37 4
721 258
721 281
644 281
644 296
5 0 17 0 0 0 0 7 0 0 37 4
548 264
548 281
544 281
544 296
5 0 17 0 0 0 0 6 0 0 37 2
435 265
435 296
0 1 17 0 0 0 0 0 8 37 0 4
644 156
644 170
721 170
721 183
0 1 17 0 0 0 0 0 7 37 0 4
544 156
544 170
548 170
548 189
1 0 17 0 0 0 0 6 0 0 37 2
435 190
435 156
0 1 17 0 0 0 0 0 5 37 0 3
327 156
329 156
329 190
1 0 17 0 0 4224 0 3 0 0 0 4
171 156
731 156
731 296
171 296
1
-21 0 0 0 700 0 0 0 0 3 2 1 34
14 Century Gothic
0 0 0 13
758 21 951 56
768 29 940 54
13 JOHN REY MOZO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
